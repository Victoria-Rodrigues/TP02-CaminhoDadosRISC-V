module add(
    input [63:0] valor1,
    input [63:0] valor2,
    output [63:0] saida
);
    assign saida = valor1 + valor2;
    
endmodule

    